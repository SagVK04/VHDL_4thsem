module new;
    initial begin
        $display("Hello World!");
    end
endmodule
